{"parameters":[{"defender":"HumanPlayer"},{"attacker":"AIRandom"},{"winner":"None"},{"playingPlayer":"Defender"},{"plays":"(4,1) (1,7))4,1()1,7(\n(4,5) (5,2))4,5()5,2(\n(3,8) (6,3))3,8()6,3(\n"}]}
{"board":"G # # AT AT AT # # G \n# # # # AT # # # # \n# # # # DT DT # # # \nAT # # # DT # AT # # \nAT # DT DT K # DT AT AT \nAT # # # DT # # # AT \n# # # # DT # # # # \n# AT # # AT # # # # \nG # # AT AT AT # # G \n"}
